module twinactions

pub struct MyStruct {
pub mut:
	a string
}

// rought splitter for json, splits a list of dicts into the text blocks
pub fn test(r string, clean bool) {

}

