module websocket

const deploy_machines_form = websocket.Form{
	q_type: websocket.q_types.form,
	question: '# Deploy a Virtual Machine',
	chat_id: "0",
	id: 10,
	description: 'VM Deployment Spces',
	form: [
		websocket.QuestionInput{
		q_type: websocket.q_types.input,
		id: id++,
		question: '### What is the name of your VM?',
		descr: 'VM Name',
		returntype: 'string',
		regex: '.*',
		regex_errormsg: '',
		min: 0,
		max: 0,
		sign: false,
		symbol: 'vm_name',
		answer: 'testvm',
		},
		websocket.QuestionInput{
		q_type: websocket.q_types.input,
		id: id++,
		question: '### Node ID',
		descr: '',
		returntype: 'string',
		regex: '.*',
		regex_errormsg: '',
		min: 0,
		max: 0,
		sign: false,
		symbol: 'node_id',
		answer: '11',
		},
		websocket.QuestionYn{
		q_type: websocket.q_types.yn,
		chat_id: "0",
		question: '### Public Ip',
		id: id++,
		symbol: 'public_ip',
		answer: false,
		},
		websocket.QuestionYn{
		q_type: websocket.q_types.yn,
		chat_id: "0",
		question: '### Planetry Ip',
		id: id++,
		symbol: 'planetry_ip',
		answer: true,
		},
		websocket.QuestionInput{
		q_type: websocket.q_types.input,
		id: id++,
		question: '### CPU Cores',
		descr: '',
		returntype: 'string',
		regex: '.*',
		regex_errormsg: '',
		min: 0,
		max: 0,
		sign: false,
		symbol: 'cpu',
		answer: 1,
		},
		websocket.QuestionInput{
		q_type: websocket.q_types.input,
		id: id++,
		question: '### Memory in MB',
		descr: '',
		returntype: 'string',
		regex: '.*',
		regex_errormsg: '',
		min: 0,
		max: 0,
		sign: false,
		symbol: 'memory',
		answer: 1024,
		},
		websocket.QuestionInput{
		q_type: websocket.q_types.input,
		id: id++,
		question: '### Root FS in GB',
		descr: '',
		returntype: 'string',
		regex: '.*',
		regex_errormsg: '',
		min: 0,
		max: 0,
		sign: false,
		symbol: 'root_fs',
		answer: 1,
		},
		websocket.QuestionInput{
		q_type: websocket.q_types.input,
		id: id++,
		question: '### Flist',
		descr: '',
		returntype: 'string',
		regex: '.*',
		regex_errormsg: '',
		min: 0,
		max: 0,
		sign: false,
		symbol: 'flist',
		answer: 'https://hub.grid.tf/tf-official-apps/threefoldtech-ubuntu-20.04.flist',
		},
		websocket.QuestionInput{
		q_type: websocket.q_types.input,
		id: id++,
		question: '### Entrypoint',
		descr: '',
		returntype: 'string',
		regex: '.*',
		regex_errormsg: '',
		min: 0,
		max: 0,
		sign: false,
		symbol: 'entrypoint',
		answer: '/init.sh',
		},
		websocket.QuestionInput{
		q_type: websocket.q_types.input,
		id: id++,
		question: '### SSH Key',
		descr: '',
		returntype: 'string',
		regex: '.*',
		regex_errormsg: '',
		min: 0,
		max: 0,
		sign: false,
		symbol: 'ssh_key',
		answer: '',
		},

	],
	symbol: "vm_specs"
	sign: false
}

const list_services_question = QuestionChoice{
  q_type: q_types.choices,
  question: "Choose a services",
  id: id++
  descr: "services"
  sorted: true
  choices: [
	Choice{
		value: "deploy_vm_form",
		title: "Deploy VM",
	},
	Choice{
		value: "ping",
		title: "Ping",
	}
  ]
  multi: false,
  sign: false,
  symbol: "service",

  answer: "",
}