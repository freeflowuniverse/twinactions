module main
import websocket as ws


fn main() {
	ws.serve()?
}
