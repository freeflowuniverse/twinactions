module websocket

// ERROR handlera
const (
	no_event = "There is no event to do this action."
	no_data = "You must provide a data."
)