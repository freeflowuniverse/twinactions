module websocket

const deploy_machines_form = websocket.Form{
	q_type: websocket.q_types.form,
	question: '# Deploy a Virtual Machine',
	chat_id: "0",
	id: 10,
	description: 'VM Deployment Spces',
	form: [
		websocket.QuestionInput{
		q_type: websocket.q_types.input,
		id: id++,
		question: '### What is the name of your VM?',
		descr: 'VM Name',
		returntype: 'string',
		regex: '.*',
		regex_errormsg: '',
		min: 0,
		max: 0,
		sign: false,
		symbol: 'vm_name',
		answer: '',
		},
		websocket.QuestionInput{
		q_type: websocket.q_types.input,
		id: id++,
		question: '### Node ID',
		descr: '',
		returntype: 'string',
		regex: '.*',
		regex_errormsg: '',
		min: 0,
		max: 0,
		sign: false,
		symbol: 'node_id',
		answer: '',
		},
		websocket.QuestionYn{
		q_type: websocket.q_types.yn,
		chat_id: "0",
		question: '### Public Ip',
		id: id++,
		symbol: 'public_ip',
		answer: '',
		},
		websocket.QuestionYn{
		q_type: websocket.q_types.yn,
		chat_id: "0",
		question: '### Planetry Ip',
		id: id++,
		symbol: 'planetry_ip',
		answer: '',
		},
		websocket.QuestionInput{
		q_type: websocket.q_types.input,
		id: id++,
		question: '### CPU Cores',
		descr: '',
		returntype: 'string',
		regex: '.*',
		regex_errormsg: '',
		min: 0,
		max: 0,
		sign: false,
		symbol: 'cpu',
		answer: '',
		},
		websocket.QuestionInput{
		q_type: websocket.q_types.input,
		id: id++,
		question: '### Memory in MB',
		descr: '',
		returntype: 'string',
		regex: '.*',
		regex_errormsg: '',
		min: 0,
		max: 0,
		sign: false,
		symbol: 'memory',
		answer: '',
		},
		websocket.QuestionInput{
		q_type: websocket.q_types.input,
		id: id++,
		question: '### Root FS in GB',
		descr: '',
		returntype: 'string',
		regex: '.*',
		regex_errormsg: '',
		min: 0,
		max: 0,
		sign: false,
		symbol: 'root_fs',
		answer: '',
		},
		websocket.QuestionInput{
		q_type: websocket.q_types.input,
		id: id++,
		question: '### Flist',
		descr: '',
		returntype: 'string',
		regex: '.*',
		regex_errormsg: '',
		min: 0,
		max: 0,
		sign: false,
		symbol: 'flist',
		answer: '',
		},
		websocket.QuestionInput{
		q_type: websocket.q_types.input,
		id: id++,
		question: '### Entrypoint',
		descr: '',
		returntype: 'string',
		regex: '.*',
		regex_errormsg: '',
		min: 0,
		max: 0,
		sign: false,
		symbol: 'entrypoint',
		answer: '',
		},
		websocket.QuestionInput{
		q_type: websocket.q_types.input,
		id: id++,
		question: '### SSH Key',
		descr: '',
		returntype: 'string',
		regex: '.*',
		regex_errormsg: '',
		min: 0,
		max: 0,
		sign: false,
		symbol: 'ssh_key',
		answer: '',
		},

	],
	symbol: "vm_specs"
	sign: false
}

const list_services_question = QuestionChoice{
  q_type: q_types.choices,
  question: "Choose a services",
  id: id++
  descr: "services"
  sorted: true
  choices: [
	Choice{
		value: "deploy_vm_form",
		title: "Deploy VM",
	},
	Choice{
		value: "ping",
		title: "Ping",
	}
  ]
  multi: false,
  sign: false,
  symbol: "service",

  answer: "",
}