module twinactions
